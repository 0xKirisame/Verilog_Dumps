module BCD_7SEG(X,F);
	
	input [3:0] X;
	output [6:0] F;
	
	assign F[0] = !X[3] && X[2] && !X[0] || !X[3] && !X[2] && !X[1] && X[0];
	
	assign F[1] = !X[3] && X[2] && !X[1] && X[0] || !X[3] && X[2] && X[1] && !X[0];
	
	assign F[2] = !X[3] && !X[2] && X[1] && !X[0];		 
	
	assign F[3] = !X[3] && !X[2] && !X[1] && X[0] || !X[3] && X[2] && !X[1] && !X[0] || !X[3] && X[2] && X[1] && X[0];
	
	assign F[4] = !X[3] && X[0] || !X[2] && !X[1] && X[0] || !X[3] && X[2] && !X[1];							   
	
	assign F[5] = !X[3] && !X[2] && X[0] || !X[3] && !X[2] && X[1] || !X[3] && X[1] && X[0];						
	
	assign F[6] = !X[3] && !X[2] && !X[1] || !X[3] && X[2] && X[1] && X[0];											 
	
endmodule